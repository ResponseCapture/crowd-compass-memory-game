<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 18.1.1, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
   viewBox="356 29.5 280 500" enable-background="new 356 29.5 280 500" xml:space="preserve">
<g>
  <g>
    <path fill="#FFFFFF" d="M581.1,35.1H415.3c-25.2,0-45.6,20.4-45.6,45.6v398.7c0,25.2,20.4,45.6,45.6,45.6h165.8
      c25.2,0,45.6-20.4,45.6-45.6V80.8C626.7,55.6,606.3,35.1,581.1,35.1z"/>
    <path fill="#00D6EE" d="M471.3,75.7h53.8c3.4,0,6.2-2.8,6.2-6.2c0-3.4-2.8-6.2-6.2-6.2h-53.8c-3.4,0-6.2,2.8-6.2,6.2
      C464.9,72.9,467.7,75.7,471.3,75.7z M471.3,67h53.8c1.4,0,2.2,1.1,2.2,2.2c0,1.4-1.1,2.2-2.2,2.2h-53.8c-1.4,0-2.2-1.1-2.2-2.2
      C468.8,68.2,469.9,67,471.3,67z"/>
    <path fill="#00D6EE" d="M498.2,477.8c-7.6,0-13.7,6.2-13.7,13.7c0,7.6,6.2,13.7,13.7,13.7c7.6,0,13.7-6.2,13.7-13.7
      C511.9,484,505.8,477.8,498.2,477.8z M498.2,501.3c-5.3,0-9.8-4.5-9.8-9.8c0-5.3,4.5-9.8,9.8-9.8s9.8,4.5,9.8,9.8
      C508,496.8,503.5,501.3,498.2,501.3z"/>
    <path fill="#651FFF" d="M549.2,354.6c-0.3,0-0.6,0-0.8-0.3L498.2,328l-50.1,26.3c-0.6,0.3-1.4,0.3-2.2-0.3c-0.6-0.6-0.8-1.1-0.8-2
      l9.5-55.7l-40.6-39.5c-0.6-0.6-0.8-1.4-0.6-2c0.3-0.8,0.8-1.1,1.7-1.4l56-8.1l24.9-50.7c0.3-0.6,1.1-1.1,1.7-1.1l0,0
      c0.8,0,1.4,0.6,1.7,1.1l24.9,50.7l56,8.1c0.8,0,1.4,0.6,1.7,1.4c0.3,0.8,0,1.4-0.6,2l-40.6,39.5l9.5,55.7c0,0.8-0.3,1.4-0.8,2
      C550,354.3,549.5,354.6,549.2,354.6z"/>
    <path fill="#00D6EE" d="M387.9,460.4h220.6V90.8H387.9V460.4z M604.3,95v361.5H391.8V95H604.3z"/>
  </g>
</g>
</svg>
