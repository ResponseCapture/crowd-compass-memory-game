<svg viewbox="0 0 20 20" width="15px" height="15px">
  <rect x="9" y="0" width="2" height="20" fill="#FFF" transform="rotate(45 10 10)"></rect>
  <rect x="9" y="0" width="2" height="20" fill="#FFF" transform="rotate(-45 10 10)"></rect>
</svg>