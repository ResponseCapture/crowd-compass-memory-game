<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 18.1.1, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
	 viewBox="0 0 1950 750" enable-background="new 0 0 1950 750" xml:space="preserve">
<g>
	<path fill="#283238" d="M1954.6,1139c-2.5,0-3.6,1.4-4.2,2.3v0h0c0,0,0,0,0,0v-2h-4.7c0.1,1.3,0,14.1,0,14.1h4.7v-7.9
		c0-0.4,0-0.8,0.2-1.1c0.3-0.8,1.1-1.7,2.4-1.7c1.7,0,2.4,1.3,2.4,3.2v7.5h4.7v-8.1C1959.9,1141,1957.6,1139,1954.6,1139z"/>
	<path fill="#283238" d="M1940.7,1132.5c-1.6,0-2.7,1.1-2.7,2.4c0,1.4,1,2.4,2.6,2.4h0c1.6,0,2.7-1.1,2.7-2.4
		C1943.3,1133.5,1942.3,1132.5,1940.7,1132.5z"/>
	<rect x="1938.4" y="1139.3" fill="#283238" width="4.7" height="14.1"/>
</g>
<path fill="#2F383E" d="M212.8,409.8c171.5-24.7,346.2-2.3,495.1,48.8c232.7,79.9,456.4,283,762.6,253.5
	c302.4-29.1,452.1-214.9,465.6-229.3V15H16.1v444.9C78.3,437.2,143.8,419.7,212.8,409.8z"/>
</svg>
