<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 18.1.1, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
   viewBox="397 183 162 192" enable-background="new 397 183 162 192" xml:space="preserve">
<g>
  <path fill="#FFFFFF" d="M481.1,221.2c-0.1,1.1-2.2,5.4-4.8,6c-1.2,0.4-2.9,1.3-3,2c0,0.2,0.2,0.8,2,1.6l1,0.4l1.4-0.1l0.2-0.9
    l1,0.3l-0.8,3.1c0.4,0.2,0.8,0.4,1.3,0.7c0.2,0.1,0.4,0.2,0.6,0.3l0.7,0.4c0.3,0.2,0.6,0.2,0.8,0.2c0.1,0,0.1,0,0.2,0
    c0.2-0.1,0.3-0.2,0.4-0.2l0.1-0.1c0.2-0.3,0.5-0.5,0.7-0.8c0.3-0.3,0.5-0.5,0.8-0.7l0.7-0.6l-0.6-0.7l-0.6-0.8l-0.3-0.4l0.8-0.7
    l0.9,1.2h0.6c4.1,0.2,7.6,3,9.3,4.7c0.1,0.1,0.3,0.3,0.4,0.4c1.2,1.2,2.6,2.1,4.2,2.6c0-1.4-0.2-2.2-0.2-2.2v-0.1l-6.2-33
    c-0.2-0.1-0.3-0.3-0.5-0.4l-0.2,4.1c0,0-1.2-3-2.2-3.4l-0.6,3.6c-1.8-3.7-4.6-4.5-4.6-4.5s-0.2,2.7-0.6,4.4l-6-5.6
    c-1.6-1.9-4.3-0.7-6,0.2l-2.5,8.4c2.5,0.1,7.3,0.8,10,3.8C480.9,216,481.5,218.3,481.1,221.2z M489.3,215.8c0.6,0,1,0.5,1,1
    c0,0.6-0.5,1-1,1c-0.6,0-1-0.5-1-1C488.2,216.3,488.7,215.8,489.3,215.8z"/>
  <path fill="#FFFFFF" d="M465.7,218.9c-1.3-0.3-2.7,0.5-3.2,1.8c-0.2,0.7-0.2,1.5,0.1,2.1c0.3,0.6,0.8,1.1,1.5,1.3L465.7,218.9z"/>
  <path fill="#FFFFFF" d="M466.3,235.9c1.5-1.5,4.4-3.9,7.9-4.5c-1.3-0.7-1.9-1.5-1.9-2.3c0.1-1.7,3.1-2.8,3.7-3l0,0
    c2-0.5,3.9-4.3,4-5.1c0.3-2.5-0.2-4.6-1.5-6.1c-2.5-2.8-7.2-3.4-9.5-3.5l-7,23.1c-0.5,1.6-0.9,3.1-1.4,4.5c2-0.3,3.9-1.3,5.3-2.8
    C466.1,236.2,466.2,236,466.3,235.9z M474.2,215.8c0.6,0,1,0.5,1,1c0,0.6-0.5,1-1,1c-0.6,0-1-0.5-1-1S473.7,215.8,474.2,215.8z"/>
  <path fill="#FFFFFF" d="M460,246l0.5-1c0-0.1-0.1,0.1-0.1,0.1c-0.2-0.3-0.3-0.6-0.5-0.9l0,0c-0.3,0-0.6,0-0.8,0
    c-1.7,0-3.3-0.4-4.5-0.6l-1.1,2.5h6.5V246z"/>
  <path fill="#FFFFFF" d="M453.4,243.5c-0.5-0.2-3.3-1-5.1-2.7c-0.6-0.6-1.1-1.2-1.4-1.8c-3.4-1.2-7.3-2.2-9.9-2.4l0,0l-0.3-0.1
    c-0.1,0-9.5-2.4-16,4.6l-0.8-0.7c6.3-6.7,15-5.3,16.7-4.9c1.7-1.6,2.8-4.8,3-5.2l2.8-16.5l0.1-0.6c0.4-1.8,0.6-2.9,0.4-3.3
    l-0.1-0.1c-0.5-0.8-1-1.6-1.5-2.4l-7.9-15.7c-0.5-1-1-1.6-1.7-1.7c-1-0.1-2.2,1-2.6,1.4l-7,7.8c-1.5,1.6-1.6,2.4-1.5,2.8
    c0.1,0.5,0.7,0.6,0.7,0.6l9.4,3c0.2-0.1,0.4-0.3,0.4-0.6c0.1-0.5-0.2-1.9-4.1-4.9l-0.5-0.4l2.9-2.6l0.7,0.8l-1.4,1.2l1.6,0.1v1.1
    H429c2.4,2,3.5,3.6,3.2,4.9c-0.1,0.9-0.9,1.4-1.3,1.5l-0.2,0.1l-6.1-1.9c-0.7,0.9-1.9,2.9-1.4,4.2c0.4,0.9,1.6,1.5,3.5,1.8
    l11.3,0.7l-22.5,13.3c-0.3,0.3-4.6,3.6-5.1,6.6c0,0.2-0.1,0.6-0.4,1.7c-2.5,10.3-3.7,16.8-3.5,19.4c0.4-0.4,0.7-0.8,1.2-1.2
    l0.7,0.8c-2.6,2.6-3.8,4.7-3.3,6.2c0.6,2,3.8,2.5,3.8,2.5h0.1l29.6,17.5L453.4,243.5L453.4,243.5z"/>
  <path fill="#FFFFFF" d="M499,225c0.4-0.6,0.6-1.3,0.5-2.1c-0.2-1.3-1.3-2.3-2.6-2.4l1,5.3C498.4,225.7,498.8,225.4,499,225z"/>
  <path fill="#FFFFFF" d="M480.7,248c0,0.9,0.6,1.7,1.7,2.4c2.2,1.4,5,1.7,7.5,0.6c0.5-0.2,0.9-0.4,1.4-0.7c2.9-1.5,5.1-3.8,6.4-6.6
    c-0.9-0.2-1.7-0.5-2.5-0.8c-0.1-0.1-0.6-0.3-1.1-0.5c-0.8-0.4-1.9-0.8-2.4-1.1c-3.5-1.8-7.4-2.8-11.4-3.1l0,0l0,0
    c-4,0.2-7.9,1.3-11.4,3.1c-0.6,0.3-1.6,0.7-2.4,1.1c-0.5,0.2-1,0.4-1.1,0.5c-1,0.5-2.2,0.8-3.3,1l-0.5,1.1c0.6,0.8,1.4,1.4,2.2,2
    c1.6,1,4.8,2.8,7.4,4c2.3,1.1,4.9,0.8,6.9-0.6c0.9-0.7,1.4-1.4,1.4-2.1c0-1-0.9-2.1-2.6-3.2l0.6-0.9c1.1,0.7,1.9,1.5,2.4,2.2
    c0.5-1.1,1.5-2.2,3-3.3l0.7,0.9C481.7,245.5,480.7,246.9,480.7,248z M481.7,240.3c-1.5-0.6-3.3,0.9-3.3,1l-0.7-0.8
    c0.1-0.1,2.3-2,4.4-1.2L481.7,240.3z"/>
  <path fill="#FFFFFF" d="M504.5,246l-1-2.1c-0.6,0-1.1,0.3-1.7,0.3c-0.5,0-1.1-0.1-1.7-0.2l-0.8,0.4l0.4,1.6H504.5z"/>
  <path fill="#FFFFFF" d="M457,254h-6.7l-3,7h8.4c-0.2-1-0.2-2-0.2-2.6s0.1-1.1,0.3-1.7L457,254z"/>
  <path fill="#FFFFFF" d="M479,272.9c14.9,0,22.4-4.9,22.5-14.5c0-0.4,0-0.6-0.3-1.4l-3-11.6c-1.5,2.5-3.6,4.5-6.3,5.9
    c-0.5,0.3-1,0.5-1.5,0.7c-1.2,0.5-2.5,0.8-3.7,0.8c-1.7,0-3.4-0.5-4.8-1.4c-0.7-0.5-1.2-1-1.6-1.5c-0.3,0.5-0.8,1-1.4,1.4
    c-2.3,1.6-5.3,1.9-8,0.7s-5.9-3-7.5-4c-0.8-0.5-1.5-1.1-2.2-1.8l-4.4,10.8c-0.2,0.4-0.3,0.9-0.3,1.3c0,1.5,0.3,5.5,3.6,8.9
    c0.1,0.1,0.2,0.2,0.3,0.3c0.2,0.2,0.4,0.5,0.6,0.5h0C464.8,271,470.9,272.9,479,272.9z"/>
  <path fill="#FFFFFF" d="M510.6,261l-3-7h-6.1l0.7,2.7c0.4,0.9,0.4,1.3,0.4,1.8s0,1.5-0.2,2.5H510.6z"/>
  <path fill="#FFFFFF" d="M499,268c-3.8,4-10.5,6-20,6c-9,0-15.6-2-19.6-6h-15.1l-3.1,7h75.3l-3.1-7H499z"/>
  <path fill="#FFFFFF" d="M482,327.5c5,2.4,13.4-0.1,13.4-0.1l0.2-0.1l-0.1-2.2H482V327.5z"/>
  <path fill="#FFFFFF" d="M461.4,328.8c-0.4,1.5-0.9,5.3,2.4,9.8c0.3,0.4,0.5,0.8,0.8,1.1c0.1,0.2,0.2,0.3,0.3,0.5
    c0.3,0.4,0.6,0.6,0.9,0.6c0.6,0.1,1.3-0.4,2.2-1.3l0.8,0.7c-1.1,1.1-2.1,1.7-3,1.6c-0.7-0.1-1.3-0.4-1.7-1.1
    c-0.1-0.2-0.2-0.3-0.3-0.5c-0.1-0.2-0.3-0.4-0.4-0.6c-0.1,3.2,0,6.5,0.3,9.7l0.1,0.6l6.2-0.2l1.2-9.1l0.3-0.1
    c1.9-0.9,2.9-7.3,3.2-11.8c-1.7,0.6-3.6,0.9-5.8,0.9C465.4,329.8,462.5,329.1,461.4,328.8z"/>
  <polygon fill="#FFFFFF" points="449.4,289 508.5,289 515.3,282 442.6,282   "/>
  <path fill="#FFFFFF" d="M550.4,251.3c0.4,0.4,0.8,0.8,1.2,1.2c0.2-2.6-1-9.2-3.5-19.4c-0.3-1-0.4-1.5-0.4-1.7
    c-0.5-3-4.8-6.3-5.1-6.6l-22.5-13.3l11.3-0.7c1.9-0.2,3.1-0.8,3.5-1.8c0.5-1.4-0.7-3.3-1.4-4.2l-6.1,1.9l-0.2-0.1
    c-0.4-0.1-1.1-0.6-1.3-1.5c-0.2-1.3,0.9-2.9,3.2-4.9h-1.3v-1.1l1.6-0.1l-1.4-1.2l0.7-0.8l2.9,2.6l-0.5,0.4c-4,2.9-4.2,4.4-4.1,4.9
    c0.1,0.3,0.3,0.5,0.4,0.6l9.4-3c0,0,0.6-0.2,0.7-0.6c0.1-0.4,0-1.2-1.5-2.8l-7-7.8c-0.4-0.5-1.6-1.6-2.6-1.5
    c-0.6,0.1-1.2,0.6-1.7,1.7l-7.9,15.7c-0.4,0.8-1,1.6-1.5,2.4l-0.1,0.1c-0.2,0.3,0,1.4,0.4,3.3l0.1,0.6l2.8,16.5
    c0.1,0.4,1.3,3.6,3,5.2c1.7-0.4,10.5-1.8,16.7,4.9l-0.8,0.7c-6.5-6.9-15.9-4.6-16-4.6l-0.3,0.1l0,0c-1.9,0.1-4.3,0.7-6.8,1.5
    c-0.4,0.9-1,1.9-2,2.8c-1.8,1.7-4.6,2.5-5.1,2.7c-0.6,0.2-1.4,0.3-2.5,0.5l14.4,34.3l29.6-17.5h0.1c0,0,3.2-0.5,3.8-2.5
    c0.5-1.5-0.7-3.7-3.3-6.2L550.4,251.3z"/>
  <polygon fill="#FFFFFF" points="463.2,304 494.6,304 501.4,297 456.4,297   "/>
  <polygon fill="#FFFFFF" points="494.6,311 463,311 462.4,318 495.1,318   "/>
  <path fill="#FFFFFF" d="M461.8,327.4c1.6,0.4,8.2,2.1,13.2,0.1V325h-13.2V327.4z"/>
  <path fill="#FFFFFF" d="M488,329.8c-2.2,0-4.2-0.3-5.9-0.9c0.3,4.4,1.4,10.8,3.2,11.7l0.2,0.1l1.2,9.1l6.2,0.2l0.1-0.6
    c0.3-3.2,0.5-6.5,0.3-9.7c-0.1,0.2-0.3,0.4-0.4,0.6s-0.2,0.3-0.3,0.5c-0.4,0.7-1,1-1.7,1.1c-0.9,0.1-2-0.5-3-1.6l0.8-0.7
    c0.8,0.9,1.6,1.3,2.2,1.3c0.3,0,0.7-0.2,0.9-0.6c0.1-0.2,0.2-0.3,0.3-0.5c0.2-0.4,0.5-0.8,0.8-1.1c3.2-4.4,2.8-8.1,2.4-9.7
    C493.8,329.3,491,329.8,488,329.8z"/>
  <path fill="#FFFFFF" d="M552.5,253.6c0.8-2.9-1.4-12.5-3.4-20.8c-0.2-0.8-0.4-1.5-0.4-1.6c-0.6-3.5-5.3-7.2-5.5-7.3l-19.5-11.5
    l7.8-0.5c2.4-0.3,3.9-1.1,4.4-2.4c0.7-1.8-0.6-3.9-1.3-5l2.6-0.8c0.4-0.1,1.2-0.5,1.4-1.3c0.3-1-0.3-2.3-1.7-3.8l-7-7.8
    c-0.1-0.1-1.7-2.1-3.6-1.8c-1,0.1-1.9,0.9-2.5,2.3l-7.9,15.7c-0.4,0.8-0.9,1.6-1.4,2.3l-0.1,0.1c-0.5,0.7-0.3,1.6,0.3,4.1l0.1,0.5
    l2.8,16.5v0.1c0,0.1,1.1,3.1,2.7,5.1c-1.6,0.2-3.4,0.6-5.3,1.2c0.1-0.3,0.2-0.5,0.2-0.6c1.2-5.4-1.2-8.3-3.3-9.9
    c-1.4-1-3-1.5-4.7-1.5c-0.5,0-1,0.1-1.5,0.2c-3,0.6-3.9,2.7-3.7,4.4c0.2,2.1,2,4.3,4.8,4.3c0.3,0,0.7,0,1-0.1l1.7-0.4l-1.5-1
    c-2.2-1.5-2.6-2.4-2.6-2.7c0-0.1,0-0.4,0.6-0.8c0.2-0.2,0.5-0.2,0.8-0.2c0.7,0,1.5,0.4,1.8,0.5c2,1.2,1.9,4.4,1.2,6.4
    c-1,2.9-3.1,4-7.2,4c-0.4,0-0.8,0-1.2,0c-0.2,0-0.3,0-0.5,0c-0.3,0-0.5-0.1-0.8-0.1c0.1-1.6-0.2-2.5-0.3-2.8l-1.8-9.4
    c1.7-0.6,2.7-2.3,2.5-4.2c-0.3-1.9-2-3.3-3.9-3.3l-2.7-14.2c1.3,2.1,1.7,4.4,1.7,4.4c1.9-5.7-0.4-10-1-10.9
    c-0.1-0.2-0.2-0.4-0.3-0.5c-1.4-2.7-3.5-4.2-5.6-5.1c-3.2-1.4-6.8-1.3-10.1,0c-8.6,3.4-8.2,9.7-8.2,9.7l-2.2,7.2h-0.1v0.5l-2.2,7.2
    c-1.9-0.4-3.9,0.7-4.5,2.5c-0.3,1-0.3,2,0.2,3c0.4,0.9,1.2,1.6,2.1,1.9l-2.4,7.8c-0.5,1.1-0.8,2.3-1.1,3.5
    c-0.3,0.8-0.5,1.6-0.8,2.3c0,0.1-0.1,0.3-0.1,0.4c0,0,0,0-0.1,0c-0.4,0-0.8,0-1.2,0c-4.1,0-6.2-1.2-7.2-4c-0.7-1.9-0.7-5.2,1.2-6.4
    c0.3-0.2,1.1-0.5,1.8-0.5c0.3,0,0.6,0.1,0.8,0.2c0.6,0.4,0.6,0.7,0.6,0.8c0,0.4-0.3,1.2-2.6,2.7l-1.5,1l1.7,0.4
    c0.3,0.1,0.7,0.1,1,0.1c2.7,0,4.5-2.2,4.8-4.3c0.2-1.7-0.7-3.8-3.7-4.4c-0.5-0.1-1-0.2-1.5-0.2c-1.7,0-3.3,0.5-4.7,1.5
    c-2.2,1.6-4.5,4.5-3.3,9.9c0,0.1,0.2,0.6,0.5,1.4c-2.8-0.9-5.9-1.7-8.2-2.1c1.6-2,2.7-4.9,2.7-5.1l2.8-16.6l0.1-0.6
    c0.5-2.5,0.7-3.4,0.3-4.1l-0.1-0.1c-0.5-0.7-1-1.5-1.4-2.3l-7.9-15.7c-0.6-1.4-1.5-2.2-2.5-2.3c-1.9-0.2-3.5,1.7-3.5,1.8l-7,7.8
    c-1.4,1.5-2,2.8-1.7,3.8c0.2,0.8,1,1.2,1.4,1.3l2.6,0.8c-0.7,1-2,3.2-1.3,5c0.5,1.3,2,2.2,4.4,2.5l7.8,0.5l-19.5,11.5l0,0
    c-0.2,0.2-5,3.8-5.5,7.3c0,0.1-0.2,0.8-0.4,1.6c-2,8.2-4.1,17.9-3.4,20.8c-1.4,1.9-1.9,3.6-1.5,5c0.8,2.4,3.9,3.1,4.6,3.2
    l29.6,17.5l-0.1,0.1l24.1,25.1l-2,23.3c-0.3,0.9-1.6,5.1,1.7,10.5c-0.2,3.8-0.1,7.6,0.3,11.3l0.2,1.6h0.2l0.2,10.3
    c0,0-1.1,0.2-7.9,9.1c-1.5,1.9,3.6,2.4,8.3,0.1c0.8-0.4,1.7-0.8,2.6-1.1c5.3-2.1,5.3-5.8,5.2-6.9c0-0.3-0.4-9.7-0.5-11.7l0,0
    l1.3-9.5c2.7-1.9,3.5-10.4,3.7-13l0.2-0.1V325h5v3.5l0.1,0.1c0.2,2.6,0.8,11.1,3.5,13l1.2,9.5l0,0c-0.1,2-0.5,11.4-0.5,11.7
    c-0.1,1.1,0,4.8,5.2,6.9c0.9,0.3,1.7,0.7,2.6,1.1c4.7,2.3,9.8,1.8,8.3-0.1c-6.8-8.9-7.9-9.1-7.9-9.1l0.2-10.3h0.2l0.2-1.6
    c0.4-3.7,0.5-7.6,0.3-11.3c2.7-4.3,2.4-8,2-9.6h0.1l0.4-0.1l-1.5-24l24.2-25.1l29.9-17.7c0.6-0.1,3.8-0.8,4.6-3.2
    C554.4,257.2,553.9,255.5,552.5,253.6z M500.1,244c0.6,0,1.2,0.2,1.7,0.2c0.6,0,1.2-0.3,1.7-0.3l1,2.1h-4.8l-0.4-1.6L500.1,244z
     M502.1,256.7l-0.7-2.7h6.1l3,7h-8.2c0.1-1,0.2-1.9,0.2-2.5C502.6,258,502.5,257.6,502.1,256.7z M460.5,267.5
    c-0.1-0.1-0.2-0.2-0.3-0.3c-3.3-3.4-3.6-7.3-3.6-8.9c0-0.4,0.1-0.9,0.3-1.3l4.4-10.8c0.6,0.7,1.3,1.3,2.2,1.8c1.7,1,4.9,2.8,7.5,4
    s5.7,0.9,8-0.7c0.6-0.4,1.1-0.9,1.4-1.4c0.4,0.5,0.9,1,1.6,1.5c1.4,1,3.1,1.4,4.8,1.4c1.2,0,2.5-0.3,3.7-0.8c0.5-0.2,1-0.4,1.5-0.7
    c2.7-1.4,4.9-3.5,6.3-5.9l3,11.6c0.3,0.8,0.3,1,0.3,1.4c-0.1,9.6-7.6,14.5-22.5,14.5c-8.1,0-14.2-1.9-18-4.9h0.1
    C460.9,268,460.7,267.6,460.5,267.5z M455.7,261h-8.4l3-7h6.7l-1.1,2.7c-0.2,0.5-0.3,1.1-0.3,1.7C455.5,259,455.5,260,455.7,261z
     M483,243.1c-1.5,1.1-2.5,2.2-3,3.3c-0.5-0.7-1.3-1.4-2.4-2.2l-0.6,0.9c1.7,1.1,2.6,2.3,2.6,3.2c0,0.7-0.5,1.4-1.4,2.1
    c-2,1.4-4.6,1.6-6.9,0.6c-2.6-1.2-5.8-3-7.4-4c-0.9-0.5-1.6-1.2-2.2-2l0.5-1.1c1.1-0.2,2.3-0.5,3.3-1c0.1-0.1,0.6-0.3,1.1-0.5
    c0.8-0.4,1.9-0.8,2.4-1.1c3.5-1.8,7.4-2.8,11.4-3.1l0,0l0,0c4,0.2,7.9,1.3,11.4,3.1c0.6,0.3,1.6,0.7,2.4,1.1c0.5,0.2,1,0.4,1.1,0.5
    c0.8,0.4,1.6,0.7,2.5,0.8c-1.3,2.8-3.6,5.1-6.4,6.6c-0.5,0.2-0.9,0.5-1.4,0.7c-2.5,1.1-5.3,0.9-7.5-0.6c-1.1-0.7-1.7-1.6-1.7-2.4
    c0-1.2,0.9-2.6,2.9-4.1L483,243.1z M499.6,222.9c0.1,0.7-0.1,1.5-0.5,2.1c-0.3,0.4-0.7,0.7-1.1,0.9l-1-5.3
    C498.2,220.6,499.4,221.6,499.6,222.9z M471.9,202c1.6-1,4.3-2.1,6-0.2l6,5.6c0.4-1.8,0.6-4.4,0.6-4.4s2.9,0.8,4.6,4.5l0.6-3.6
    c1,0.3,2.2,3.4,2.2,3.4l0.2-4.1c0.2,0.1,0.3,0.3,0.5,0.4l6.2,33v0.1c0,0,0.3,0.8,0.2,2.2c-1.6-0.5-3-1.3-4.2-2.6
    c-0.1-0.1-0.3-0.3-0.4-0.4c-1.7-1.7-5.1-4.5-9.3-4.7h-0.6l-0.9-1.2l-0.8,0.7l0.3,0.4l0.6,0.8l0.6,0.7l-0.7,0.6
    c-0.3,0.2-0.5,0.5-0.8,0.7c-0.3,0.3-0.5,0.5-0.7,0.8l-0.1,0.1c-0.1,0.1-0.2,0.2-0.4,0.2c-0.1,0-0.1,0-0.2,0c-0.2,0-0.4,0-0.8-0.2
    l-0.7-0.4c-0.2-0.1-0.4-0.2-0.6-0.3c-0.4-0.2-0.8-0.4-1.3-0.7l0.8-3.1l-1-0.3l-0.2,0.9l-1.4,0.1l-1-0.4c-1.8-0.8-2-1.4-2-1.6
    c0-0.7,1.8-1.6,3-2c2.6-0.6,4.6-4.9,4.8-6c0.4-2.8-0.2-5.2-1.8-7c-2.7-3-7.4-3.7-10-3.8L471.9,202z M462.6,222.8
    c-0.3-0.7-0.4-1.4-0.1-2.1c0.5-1.3,1.8-2.1,3.2-1.8l-1.6,5.3C463.4,223.9,462.9,223.4,462.6,222.8z M462,234.6l7-23.1
    c2.3,0.1,7,0.6,9.5,3.5c1.4,1.5,1.9,3.6,1.5,6.1c-0.1,0.8-1.9,4.7-4,5.1l0,0c-0.6,0.2-3.6,1.2-3.7,3c0,0.8,0.6,1.6,1.9,2.3
    c-3.5,0.6-6.4,3-7.9,4.5c-0.1,0.1-0.3,0.3-0.4,0.4c-1.4,1.5-3.3,2.5-5.3,2.8C461.1,237.7,461.6,236.2,462,234.6z M459,244.2
    c0.3,0,0.6,0,0.8,0l0,0c0.1,0.3,0.3,0.6,0.5,0.9c0,0.1,0.1-0.1,0.1-0.1l-0.5,1h-6.5l1.1-2.5C455.7,243.8,457.3,244.2,459,244.2z
     M409.2,260.8h-0.1c0,0-3.2-0.5-3.8-2.5c-0.5-1.5,0.6-3.7,3.3-6.2l-0.7-0.8c-0.4,0.4-0.8,0.8-1.2,1.2c-0.2-2.6,1-9.2,3.5-19.4
    c0.3-1,0.4-1.5,0.4-1.7c0.5-3,4.8-6.3,5.1-6.6l22.5-13.3l-11.3-0.7c-2-0.2-3.1-0.8-3.5-1.8c-0.5-1.4,0.7-3.3,1.4-4.2l6.1,1.9
    l0.2-0.1c0.4-0.1,1.1-0.6,1.3-1.5c0.2-1.3-0.9-2.9-3.2-4.9h1.3v-1.1l-1.6-0.1l1.4-1.2l-0.7-0.8l-2.9,2.6l0.5,0.4
    c3.9,2.9,4.2,4.4,4.1,4.9c0,0.3-0.3,0.5-0.4,0.6l-9.4-3c0,0-0.5-0.2-0.7-0.6c-0.1-0.4,0-1.2,1.5-2.8l7-7.8c0.4-0.4,1.5-1.6,2.6-1.4
    c0.6,0.1,1.2,0.6,1.7,1.7l7.9,15.7c0.4,0.8,1,1.6,1.5,2.4l0.1,0.1c0.2,0.3,0,1.4-0.4,3.3l-0.1,0.6l-2.8,16.5
    c-0.1,0.4-1.3,3.6-3,5.2c-1.7-0.4-10.5-1.8-16.7,4.9l0.8,0.7c6.5-6.9,15.9-4.6,16-4.6l0.3,0.1l0,0c2.6,0.2,6.5,1.3,9.9,2.4
    c0.4,0.6,0.8,1.3,1.4,1.8c1.8,1.7,4.6,2.5,5.1,2.7h0.1l-14.6,34.8L409.2,260.8z M471.3,340.7l-0.3,0.1l-1.2,9.1l-6.2,0.2l-0.1-0.6
    c-0.3-3.2-0.5-6.5-0.3-9.7c0.1,0.2,0.3,0.4,0.4,0.6s0.2,0.3,0.3,0.5c0.4,0.7,1,1,1.7,1.1c0.9,0.1,2-0.5,3-1.6l-0.8-0.7
    c-0.8,0.9-1.6,1.3-2.2,1.3c-0.3,0-0.7-0.2-0.9-0.6c-0.1-0.2-0.2-0.3-0.3-0.5c-0.2-0.4-0.5-0.8-0.8-1.1c-3.3-4.6-2.8-8.4-2.4-9.8
    c1.1,0.3,4.1,1,7.4,1c2.2,0,4.1-0.3,5.8-0.9C474.2,333.4,473.2,339.7,471.3,340.7z M475,327.5c-5,2-11.6,0.4-13.2-0.1V325H475
    V327.5z M462.4,318l0.6-7h31.6l0.4,7H462.4z M492.8,338.7c-0.3,0.4-0.5,0.8-0.8,1.1c-0.1,0.2-0.2,0.3-0.3,0.5
    c-0.3,0.4-0.6,0.6-0.9,0.6c-0.6,0.1-1.3-0.4-2.2-1.3l-0.8,0.7c1.1,1.1,2.1,1.7,3,1.6c0.7-0.1,1.3-0.4,1.7-1.1
    c0.1-0.2,0.2-0.3,0.3-0.5c0.1-0.2,0.3-0.4,0.4-0.6c0.1,3.2,0,6.5-0.3,9.7l-0.1,0.6l-6.2-0.2l-1.2-9.1l-0.2-0.1
    c-1.9-0.9-2.9-7.3-3.2-11.7c1.7,0.6,3.7,0.9,5.9,0.9c3.1,0,5.8-0.5,7.3-0.9C495.7,330.5,496,334.2,492.8,338.7z M495.5,325l0.1,2.2
    l-0.2,0.1c-0.1,0-8.4,2.5-13.4,0.1V325H495.5z M494.6,304h-31.4l-6.8-7h45L494.6,304z M508.5,289h-59l-6.8-7h72.7L508.5,289z
     M441.3,275l3.1-7h15.1c4,4,10.5,6,19.6,6c9.5,0,16.2-2,20-6h14.5l3.1,7H441.3z M552.9,258.3c-0.6,2-3.8,2.5-3.8,2.5H549
    l-29.6,17.5L505,244c1-0.1,1.9-0.3,2.5-0.5c0.5-0.2,3.3-1,5.1-2.7c0.9-0.9,1.5-1.9,2-2.8c2.5-0.7,4.9-1.3,6.8-1.5l0,0l0.3-0.1
    c0.1,0,9.5-2.4,16,4.6l0.8-0.7c-6.3-6.7-15-5.3-16.7-4.9c-1.7-1.6-2.8-4.8-3-5.2l-2.8-16.5l-0.1-0.6c-0.4-1.8-0.6-2.9-0.4-3.3
    l0.1-0.1c0.5-0.8,1-1.6,1.5-2.4l7.9-15.7c0.5-1,1-1.6,1.7-1.7c1-0.1,2.2,1,2.6,1.5l7,7.8c1.5,1.6,1.6,2.4,1.5,2.8
    c-0.1,0.5-0.7,0.6-0.7,0.6l-9.4,3c-0.1-0.1-0.4-0.3-0.4-0.6c-0.1-0.5,0.2-1.9,4.1-4.9l0.5-0.4l-2.9-2.6l-0.7,0.8l1.4,1.2l-1.6,0.1
    v1.1h1.3c-2.4,2-3.5,3.6-3.2,4.9c0.1,0.9,0.9,1.4,1.3,1.5l0.2,0.1l6.1-1.9c0.7,0.9,1.9,2.9,1.4,4.2c-0.4,0.9-1.6,1.5-3.5,1.8
    l-11.3,0.7l22.5,13.3c0.3,0.3,4.6,3.6,5.1,6.6c0,0.2,0.1,0.6,0.4,1.7c2.5,10.3,3.7,16.8,3.5,19.4c-0.4-0.4-0.7-0.8-1.2-1.2
    l-0.7,0.8C552.3,254.6,553.4,256.8,552.9,258.3z"/>
  <path fill="#FFFFFF" d="M477.6,240.5l0.7,0.8c0,0,1.8-1.6,3.3-1l0.4-1C479.9,238.5,477.7,240.4,477.6,240.5z"/>
  <circle fill="#FFFFFF" cx="474.2" cy="216.8" r="1"/>
  <circle fill="#FFFFFF" cx="489.3" cy="216.8" r="1"/>
</g>
<g>
  <g>
    <g>
      <path fill="#00B8D4" d="M474.2,230.6c-0.4-0.4-0.8-0.7-1.1-1.1C473.3,229.8,473.7,230.2,474.2,230.6z"/>
    </g>
    <g>
      <polygon fill="#00B8D4" points="479,322.2 475.7,322.2 475.7,325.2 481.9,325.2 481.9,322.2       "/>
    </g>
    <g>
      <path fill="#00B8D4" d="M459.9,239.7l2.7-9C461,233.1,460.1,236.4,459.9,239.7z"/>
    </g>
    <g>
      <g>
        <g>
          <g>
            <path fill="#00B8D4" d="M439.3,279.8l-30.5-18c-0.6-0.1-3.8-0.8-4.6-3.2c-0.6-2,0.6-4.4,3.6-7.3l0.7,0.8
              c-2.6,2.6-3.8,4.7-3.3,6.2c0.6,2,3.8,2.5,3.8,2.5h0.1l29.6,17.5l15.4-36.6c-2.4-0.9-12.4-4.9-17.5-5.2l0.1-1.1
              c5.9,0.4,17.8,5.3,18.3,5.5l0.5,0.2L439.3,279.8z"/>
          </g>
          <g>
            <path fill="#00B8D4" d="M405.9,253.9c-1-2.4,1.2-12.6,3.3-21.1c0.2-0.8,0.4-1.5,0.4-1.6c0.6-3.5,5.3-7.2,5.5-7.3l0,0
              l19.5-11.5l-7.8-0.5c-2.4-0.3-3.9-1.1-4.4-2.5c-0.9-2.4,1.7-5.5,1.8-5.6l0.8,0.7c-0.6,0.7-2.2,3-1.6,4.5
              c0.4,0.9,1.6,1.5,3.5,1.8l11.3,0.7l-22.5,13.3c-0.3,0.3-4.6,3.6-5.1,6.6c0,0.2-0.1,0.6-0.4,1.7c-2.9,11.9-4,18.8-3.3,20.4
              L405.9,253.9z"/>
          </g>
          <g>
            <path fill="#00B8D4" d="M420.6,241.1l-0.8-0.7c6.3-6.7,15-5.3,16.7-4.9c1.7-1.6,2.8-4.8,3-5.2l2.8-16.5l0.1-0.6
              c0.4-1.8,0.6-2.9,0.4-3.3l-0.1-0.1c-0.5-0.8-1-1.6-1.5-2.4l-7.9-15.7c-0.5-1-1-1.6-1.7-1.7c-1-0.1-2.2,1-2.6,1.4l-7,7.8
              c-1.5,1.6-1.6,2.4-1.5,2.8c0.1,0.5,0.7,0.6,0.7,0.6l9.4,3c0.2-0.1,0.4-0.3,0.4-0.6c0.1-0.5-0.2-1.9-4.1-4.9l-0.5-0.4l2.9-2.6
              l0.7,0.8l-1.9,1.7c2.9,2.3,4.3,4.1,4,5.5c-0.1,0.9-0.9,1.4-1.3,1.5l-0.2,0.1l-9.8-3.1c-0.4-0.1-1.2-0.5-1.4-1.3
              c-0.3-1,0.3-2.3,1.7-3.8l7-7.8c0.1-0.1,1.7-2,3.5-1.8c1,0.1,1.9,0.9,2.5,2.3l7.9,15.7c0.4,0.8,0.9,1.6,1.4,2.3l0.1,0.1
              c0.5,0.7,0.3,1.6-0.3,4.1l-0.1,0.6l-2.8,16.6c-0.1,0.2-1.4,4-3.5,5.9l-0.2,0.2l-0.3-0.1C436.5,236.5,427.1,234.1,420.6,241.1z
              "/>
          </g>
          <g>
            
              <rect x="427.4" y="199.3" transform="matrix(-0.9994 -3.443791e-02 3.443791e-02 -0.9994 850.656 414.3491)" fill="#00B8D4" width="3" height="1.1"/>
          </g>
          <g>
            <path fill="#00B8D4" d="M518.9,279.8l-16.3-38.7l0.5-0.2c0.5-0.2,12.4-5.1,18.3-5.5l0.1,1.1c-5.1,0.3-15.1,4.2-17.5,5.2
              l15.4,36.6l29.6-17.5h0.1c0,0,3.2-0.5,3.8-2.5c0.5-1.5-0.7-3.7-3.3-6.2l0.7-0.8c3,2.9,4.2,5.4,3.6,7.3
              c-0.8,2.4-3.9,3.1-4.6,3.2L518.9,279.8z"/>
          </g>
          <g>
            <path fill="#00B8D4" d="M552.4,253.9l-1-0.4c0.7-1.6-0.4-8.5-3.3-20.4c-0.3-1-0.4-1.5-0.4-1.7c-0.5-3-4.8-6.3-5.1-6.6
              l-22.5-13.3l11.3-0.7c1.9-0.2,3.1-0.8,3.5-1.8c0.6-1.5-1-3.8-1.6-4.5l0.8-0.7c0.1,0.1,2.7,3.2,1.8,5.6c-0.5,1.3-2,2.2-4.4,2.4
              l-7.8,0.5l19.5,11.5c0.2,0.2,5,3.8,5.5,7.3c0,0.1,0.2,0.8,0.4,1.6C551.2,241.4,553.4,251.5,552.4,253.9z"/>
          </g>
          <g>
            <path fill="#00B8D4" d="M537.6,241.1c-6.5-6.9-15.9-4.6-16-4.6l-0.3,0.1l-0.2-0.2c-2.1-1.9-3.4-5.7-3.5-5.9v-0.1l-2.8-16.5
              l-0.1-0.5c-0.5-2.5-0.7-3.4-0.3-4.1l0.1-0.1c0.5-0.7,1-1.5,1.4-2.3l7.9-15.7c0.6-1.4,1.5-2.1,2.5-2.3c1.9-0.2,3.5,1.7,3.6,1.8
              l7,7.8c1.4,1.5,2,2.8,1.7,3.8c-0.2,0.8-1,1.2-1.4,1.3l-9.7,3.1l-0.2-0.1c-0.4-0.1-1.1-0.6-1.3-1.5c-0.2-1.4,1.1-3.2,4-5.5
              l-1.9-1.7l0.7-0.8l2.9,2.6l-0.5,0.4c-4,2.9-4.2,4.4-4.1,4.9c0.1,0.3,0.3,0.5,0.4,0.6l9.4-3c0,0,0.6-0.2,0.7-0.6
              c0.1-0.4,0-1.2-1.5-2.8l-7-7.8c-0.4-0.5-1.6-1.6-2.6-1.5c-0.6,0.1-1.2,0.6-1.7,1.7l-7.9,15.7c-0.4,0.8-1,1.6-1.5,2.4l-0.1,0.1
              c-0.2,0.3,0,1.4,0.4,3.3l0.1,0.6l2.8,16.5c0.1,0.4,1.3,3.6,3,5.2c1.7-0.4,10.5-1.8,16.7,4.9L537.6,241.1z"/>
          </g>
          <g>
            
              <rect x="528.7" y="198.3" transform="matrix(-3.450166e-02 -0.9994 0.9994 -3.450166e-02 347.816 735.6899)" fill="#00B8D4" width="1.1" height="3"/>
          </g>
        </g>
        <g>
          <g>
            <polygon fill="#00B8D4" points="455.9,296.7 502,296.7 508.9,289.4 449,289.4             "/>
          </g>
          <g>
            <polygon fill="#00B8D4" points="461.5,325.2 475.7,325.2 475.7,322.6 479,322.6 481.7,322.6 481.7,325.2 496.3,325.2 
              495.8,318.1 462.1,318.1             "/>
          </g>
          <g>
            <polygon fill="#00B8D4" points="463.2,304.1 462.6,310.8 495.3,310.8 494.8,304.1 495.1,303.8 462.8,303.8             "/>
          </g>
          <g>
            <polygon fill="#00B8D4" points="508.2,253.8 505.2,246.5 498.9,246.5 500.5,253.8             "/>
          </g>
          <g>
            <path fill="#00B8D4" d="M497.5,267.9h16.7l-3-7.1h-9.4C501.5,263,500.4,265.8,497.5,267.9z"/>
          </g>
          <g>
            <polygon fill="#00B8D4" points="517.3,275.2 440.7,275.2 439.1,279.1 442.2,282.3 515.8,282.3 518.9,279.1             "/>
          </g>
          <g>
            <path fill="#00B8D4" d="M456.4,260.9h-9.7l-3,7.1h17.4C458.2,265.8,456.9,263,456.4,260.9z"/>
          </g>
          <g>
            <polygon fill="#00B8D4" points="460.4,246.5 452.8,246.5 449.7,253.8 457.5,253.8             "/>
          </g>
        </g>
      </g>
      <g>
        <path fill="#00B8D4" d="M488,329.8c-2.7,0-5-0.4-6.9-1.2l-0.3-0.1v-4.8h-5v4.8l-0.3,0.1c-1.9,0.8-4.1,1.2-6.7,1.2
          c-4.2,0-7.8-1.1-7.9-1.2l-0.4-0.1l2-24l-24.1-25.1l16.2-38.4l7.6,2.9l-5.3,13.1c-0.2,0.4-0.3,0.9-0.3,1.3c0,1.5,0.3,5.5,3.6,8.9
          c3.7,3.8,10.1,5.7,18.8,5.7c14.9,0,22.4-4.9,22.5-14.5c0-0.4,0-0.6-0.3-1.4l-3.3-13l5.5-3.1l16.2,38.5l-24.2,25.1l1.5,24
          l-0.4,0.1C496.2,328.7,492.4,329.8,488,329.8z M481.9,327.8c1.7,0.7,3.7,1,6.1,1c3.4,0,6.6-0.7,7.7-1l-1.4-23.6l0.2-0.2
          l23.9-24.8l-15.5-36.8l-3.5,2.3l2.9,12c0.4,0.9,0.4,1.3,0.4,1.8c0,1.5,0,5.6-3.2,9.2c-3.7,4.2-10.6,6.4-20.4,6.4
          c-9.1,0-15.7-2-19.6-6c-3.6-3.7-3.9-8-3.9-9.6c0-0.6,0.1-1.1,0.3-1.7l4.9-12.1l-5.6-2.1l-15.6,36.8l24,24.9l-2,23.6
          c1,0.3,3.9,1,7.2,1c2.3,0,4.2-0.3,5.9-1v-5.2h7.1v5.1H481.9z"/>
      </g>
    </g>
    <path fill="#00B8D4" d="M496,327.7l-0.2-0.4l-0.5,0.1c-0.1,0-8.1,2.5-13.7,0l-0.8-0.3v0.9c0.1,1.2,0.6,11.5,3.6,13.6l1.3,9.5
      l8.1,0.3l0.2-1.6c0.4-3.7,0.5-7.6,0.3-11.3C498.1,332.5,496.1,327.9,496,327.7z M493,349.5l-0.1,0.6l-6.2-0.2l-1.2-9.1l-0.3-0.1
      c-1.9-1-2.9-7.5-3.2-12c5.1,1.8,11.3,0.4,13.1-0.1c0.4,1.3,1.1,5.3-2.3,10.1c-0.3,0.4-0.5,0.8-0.8,1.1c-0.1,0.2-0.2,0.3-0.3,0.5
      c-0.3,0.4-0.6,0.6-0.9,0.6c-0.6,0.1-1.3-0.4-2.2-1.3l-0.8,0.7c1.1,1.1,2.1,1.7,3,1.6c0.7-0.1,1.3-0.4,1.7-1.1
      c0.1-0.2,0.2-0.3,0.3-0.5c0.1-0.2,0.3-0.4,0.4-0.6C493.5,343,493.4,346.3,493,349.5z"/>
    <path fill="#00B8D4" d="M501.4,370.7c-6.8-8.9-7.9-9.1-7.9-9.1l0.2-11.2l-7.9,0.1c0,0-0.5,11.9-0.5,12.2c-0.1,1.1,0,4.8,5.2,6.9
      c0.9,0.3,1.7,0.7,2.6,1.1C497.8,373,502.9,372.6,501.4,370.7z"/>
    <path fill="#00B8D4" d="M474.9,327.4c-5.6,2.5-13.6,0-13.7,0l-0.5-0.1l-0.2,0.4c-0.1,0.2-2,4.8,1.7,10.6
      c-0.2,3.8-0.1,7.6,0.3,11.3l0.2,1.6l8.1-0.3l1.3-9.5c3-2.1,3.6-12.4,3.6-13.6v-0.9L474.9,327.4z M471.1,340.8l-1.2,9.1l-6.2,0.2
      l-0.1-0.6c-0.3-3.2-0.5-6.5-0.3-9.7c0.1,0.2,0.3,0.4,0.4,0.6s0.2,0.3,0.3,0.5c0.4,0.7,1,1,1.7,1.1c0.9,0.1,2-0.5,3-1.6l-0.8-0.7
      c-0.8,0.9-1.6,1.3-2.2,1.3c-0.3,0-0.7-0.2-0.9-0.6c-0.1-0.2-0.2-0.3-0.3-0.5c-0.2-0.4-0.5-0.8-0.8-1.1c-3.5-4.8-2.7-8.8-2.3-10.1
      c1.8,0.5,8.1,1.9,13.1,0.1c-0.3,4.5-1.3,11-3.2,12L471.1,340.8z"/>
    <path fill="#00B8D4" d="M471.3,362.7c0-0.3-0.5-12.2-0.5-12.2l-7.9-0.1l0.2,11.2c0,0-1.1,0.2-7.9,9.1c-1.5,1.9,3.6,2.4,8.3,0.1
      c0.8-0.4,1.7-0.8,2.6-1.1C471.3,367.6,471.4,363.8,471.3,362.7z"/>
    <g>
      <g>
        <path fill="#00B8D4" d="M463.9,225.2c-1-0.3-1.8-1-2.2-1.9c-0.4-0.9-0.5-2-0.2-2.9c0.7-2,2.9-3.1,4.9-2.4l-0.3,1
          c-1.4-0.5-3,0.3-3.5,1.7c-0.2,0.7-0.2,1.5,0.1,2.1c0.3,0.7,0.9,1.2,1.6,1.4L463.9,225.2z"/>
      </g>
    </g>
    <g>
      <g>
        <path fill="#00B8D4" d="M497.4,227.1l-0.2-1.1c0.7-0.1,1.4-0.5,1.8-1.1s0.6-1.3,0.5-2.1c-0.2-1.5-1.6-2.6-3.1-2.4l-0.2-1.1
          c2.1-0.3,4,1.2,4.3,3.3C500.9,224.9,499.5,226.8,497.4,227.1z"/>
      </g>
    </g>
    <g>
      <path fill="#00B8D4" d="M486.7,252.8c-1.7,0-3.4-0.5-4.8-1.4c-0.7-0.5-1.2-1-1.6-1.5c-0.3,0.5-0.8,1-1.4,1.4
        c-2.3,1.6-5.3,1.9-8,0.7s-5.9-3-7.5-4c-1.3-0.7-2.3-1.7-3-2.9c-1.7-2.7-1.2-5-0.8-6.2c0.5-1.5,1-2.9,1.5-4.5l10.5-34.6H493
        l6.9,36.7c0.1,0.4,0.8,2.6-0.4,6.1c-1.2,3.8-3.9,6.9-7.6,8.8c-0.5,0.3-1,0.5-1.5,0.7C489.2,252.5,488,252.8,486.7,252.8z
         M483,243.1l0.7,0.9c-2,1.5-3,2.9-2.9,4.1c0,0.9,0.6,1.7,1.7,2.4c2.2,1.4,5,1.7,7.5,0.6c0.5-0.2,0.9-0.4,1.4-0.7
        c3.4-1.8,6-4.7,7.1-8.2c1.1-3.4,0.4-5.5,0.4-5.5v-0.1l-6.7-35.8h-19.8L462,234.6c-0.5,1.6-0.9,3.1-1.5,4.6c-0.3,1-0.7,3,0.7,5.3
        c0.6,1,1.6,1.9,2.7,2.6c1.6,1,4.8,2.8,7.4,4c2.3,1.1,4.9,0.8,6.9-0.6c0.9-0.7,1.4-1.4,1.4-2.1c0-1-0.9-2.1-2.6-3.2l0.6-0.9
        c1.1,0.7,1.9,1.5,2.4,2.2C480.5,245.3,481.5,244.2,483,243.1z"/>
    </g>
    <g>
      <path fill="#00B8D4" d="M478.3,241.3l-0.7-0.8c0.1-0.1,2.3-2,4.4-1.2l-0.4,1C480.1,239.7,478.4,241.3,478.3,241.3z"/>
    </g>
    <g>
      <circle fill="#00B8D4" cx="474.2" cy="216.8" r="1"/>
    </g>
    <g>
      <path fill="#00B8D4" d="M477.7,233l-2.8-1.2c-1.8-0.8-2.7-1.7-2.6-2.7c0.1-1.7,3.1-2.8,3.7-3l0,0c2-0.5,3.9-4.3,4-5.1
        c0.3-2.5-0.2-4.6-1.5-6.1c-2.9-3.3-8.7-3.5-10.4-3.5v-1.1c1.8,0,8,0.2,11.2,3.8c1.6,1.8,2.2,4.1,1.8,7c-0.2,1.1-2.2,5.4-4.8,6
        c-1.2,0.4-2.9,1.3-3,2c0,0.2,0.2,0.8,2,1.6l2.8,1.2L477.7,233z"/>
    </g>
    <g>
      <path fill="#00B8D4" d="M489.2,207.5l0.6-3.6c1,0.3,2.2,3.4,2.2,3.4l0.2-4.1c2.9,2,3.6,6.5,3.6,6.5c1.9-5.7-0.4-10-1-10.9
        c-0.1-0.2-0.2-0.4-0.3-0.5c-1.4-2.7-3.5-4.2-5.6-5.1c-3.2-1.4-6.8-1.3-10.1,0c-8.6,3.4-8.2,9.9-8.2,9.9s4.9-4,7.4-1.2l6,5.6
        c0.4-1.8,0.6-4.4,0.6-4.4S487.4,203.8,489.2,207.5z"/>
    </g>
    <g>
      <circle fill="#00B8D4" cx="489.3" cy="216.8" r="1"/>
    </g>
    <path fill="#00B8D4" d="M511.8,226.3c-1.4-1-3-1.5-4.7-1.5c-0.5,0-1,0.1-1.5,0.2c-3,0.6-3.9,2.7-3.7,4.4c0.2,2.1,2,4.3,4.8,4.3
      c0.3,0,0.7,0,1-0.1l1.7-0.4l-1.5-1c-2.2-1.5-2.6-2.4-2.6-2.7c0-0.1,0-0.4,0.6-0.8c0.2-0.2,0.5-0.2,0.8-0.2c0.7,0,1.5,0.4,1.8,0.5
      c2,1.2,1.9,4.4,1.2,6.4c-1,2.9-3.1,4-7.2,4c-0.4,0-0.8,0-1.2,0c-0.2,0-0.3,0-0.5,0c-2.3-0.2-4.5-1.2-6.1-2.9
      c-0.1-0.1-0.3-0.3-0.4-0.4c-1.7-1.7-5.1-4.5-9.3-4.7h-0.6l-0.9-1.2l-0.8,0.7l0.3,0.4l0,0l0.6,0.8l0.6,0.7l-0.7,0.6
      c-0.3,0.2-0.5,0.5-0.8,0.7c-0.3,0.3-0.5,0.5-0.7,0.8l-0.1,0.1c-0.1,0.1-0.2,0.2-0.4,0.2c-0.1,0-0.1,0-0.2,0c-0.2,0-0.4,0-0.8-0.2
      l-0.7-0.4c-0.2-0.1-0.4-0.2-0.6-0.3c-0.4-0.2-0.8-0.4-1.3-0.7l0.8-3.1l-1-0.3l-0.2,0.9l-2.2,0.1c-4.1,0.2-7.6,3-9.3,4.7
      c-0.1,0.1-0.3,0.3-0.4,0.4c-1.6,1.7-3.8,2.7-6.1,2.9c-0.1,0-0.3,0-0.5,0c-0.4,0-0.8,0-1.2,0c-4.1,0-6.2-1.2-7.2-4
      c-0.7-1.9-0.7-5.2,1.2-6.4c0.3-0.2,1.1-0.5,1.8-0.5c0.3,0,0.6,0.1,0.8,0.2c0.6,0.4,0.6,0.7,0.6,0.8c0,0.4-0.3,1.2-2.6,2.7l-1.5,1
      l1.7,0.4c0.3,0.1,0.7,0.1,1,0.1c2.7,0,4.5-2.2,4.8-4.3c0.2-1.7-0.7-3.8-3.7-4.4c-0.5-0.1-1-0.2-1.5-0.2c-1.7,0-3.3,0.5-4.7,1.5
      c-2.2,1.6-4.5,4.5-3.3,9.9c0,0.1,0.7,2.8,2.6,4.6c1.8,1.7,4.6,2.5,5.1,2.7c1.1,0.3,3.3,0.7,5.7,0.7l0,0c1.8,0,4.4-0.2,6.4-1.2
      c0.1-0.1,0.6-0.3,1.1-0.5c0.8-0.4,1.9-0.8,2.4-1.1c3.5-1.8,7.4-2.8,11.4-3.1l0,0l0,0c4,0.2,7.9,1.3,11.4,3.1
      c0.6,0.3,1.6,0.7,2.4,1.1c0.5,0.2,1,0.4,1.1,0.5c2,1,4.6,1.2,6.4,1.2c2.4,0,4.6-0.3,5.7-0.7c0.5-0.2,3.3-1,5.1-2.7
      c1.9-1.8,2.6-4.5,2.6-4.6C516.4,230.8,514,227.8,511.8,226.3z"/>
  </g>
</g>
</svg>
