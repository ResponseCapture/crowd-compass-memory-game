<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 18.1.1, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
	 viewBox="0 0 25 25" enable-background="new 0 0 25 25" xml:space="preserve">
<path fill="#283238" d="M18.2,8.2h-3.5V5.9c0-0.9,0.6-1.1,1-1.1c0.4,0,2.5,0,2.5,0V1.1l-3.4,0c-3.8,0-4.6,2.8-4.6,4.6v2.5H8v3.9h2.2
	c0,5,0,11,0,11h4.6c0,0,0-6.1,0-11h3.1L18.2,8.2z"/>
</svg>
