<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 18.1.1, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
	 viewBox="0 0 1950 500" enable-background="new 0 0 1950 500" xml:space="preserve">
<g>
	<path fill="#283238" d="M1954.6,1014c-2.5,0-3.6,1.4-4.2,2.3v0h0c0,0,0,0,0,0v-2h-4.7c0.1,1.3,0,14.1,0,14.1h4.7v-7.9
		c0-0.4,0-0.8,0.2-1.1c0.3-0.8,1.1-1.7,2.4-1.7c1.7,0,2.4,1.3,2.4,3.2v7.5h4.7v-8.1C1959.9,1016,1957.6,1014,1954.6,1014z"/>
	<path fill="#283238" d="M1940.7,1007.5c-1.6,0-2.7,1.1-2.7,2.4c0,1.4,1,2.4,2.6,2.4h0c1.6,0,2.7-1.1,2.7-2.4
		C1943.3,1008.5,1942.3,1007.5,1940.7,1007.5z"/>
	<rect x="1938.4" y="1014.3" fill="#283238" width="4.7" height="14.1"/>
</g>
<path fill="#353E44" d="M284.8,246.1c243.1,27.8,401.9,177.7,650.6,199.2c253.4,21.9,521.8-30.4,736-106
	c103-36.3,256.7-118.5,265.6-122.9V38H17v259.6C92.3,259.9,180.2,234.1,284.8,246.1z"/>
</svg>
