<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 18.1.1, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
	 viewBox="120 1 720 558" enable-background="new 120 1 720 558" xml:space="preserve">
<rect x="120.7" y="1" fill="#00E676" width="719.3" height="557.1"/>
<path opacity="0.65" fill="#69F0AE" enable-background="new    " d="M765.7,416c-64.3,8.8-129.6,0.9-185.6-17.7
	c-87.1-28.8-170.9-102.5-285.7-91.8c-113.3,10.5-169.3,77.9-174.4,83V559h719.3V397.9C816.1,406,791.7,412.5,765.7,416z"/>
</svg>
