<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 18.1.1, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
	 viewBox="0 0 600 600" enable-background="new 0 0 600 600" xml:space="preserve">
<g>
	<path fill="#283238" d="M1279.6,1064c-2.5,0-3.6,1.4-4.2,2.3v0h0c0,0,0,0,0,0v-2h-4.7c0.1,1.3,0,14.1,0,14.1h4.7v-7.9
		c0-0.4,0-0.8,0.2-1.1c0.3-0.8,1.1-1.7,2.4-1.7c1.7,0,2.4,1.3,2.4,3.2v7.5h4.7v-8.1C1284.9,1066,1282.6,1064,1279.6,1064z"/>
	<path fill="#283238" d="M1265.7,1057.5c-1.6,0-2.7,1.1-2.7,2.4c0,1.4,1,2.4,2.6,2.4h0c1.6,0,2.7-1.1,2.7-2.4
		C1268.3,1058.5,1267.3,1057.5,1265.7,1057.5z"/>
	<rect x="1263.4" y="1064.3" fill="#283238" width="4.7" height="14.1"/>
</g>
<g>
	<path fill="#7C4DFF" d="M27.5,27.6c-0.5,0-1,0.4-1,1v548c0,0.6,0.5,1,1,1h548c0.5,0,1-0.4,1-1v-548c0-0.6-0.5-1-1-1H27.5z
		 M565.5,565.6c0,0.6-0.5,1-1,1h-526c-0.6,0-1-0.4-1-1v-526c0-0.5,0.4-1,1-1h526c0.5,0,1,0.5,1,1V565.6z"/>
</g>
</svg>
