<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 18.1.1, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
	 viewBox="576.3 239.6 605 550" enable-background="new 576.3 239.6 605 550" xml:space="preserve">
<path fill="#F1F4F5" d="M1170.7,400.7c-2.2-172.1-220.5-220.9-294.2-58.4c-76.7-161.2-295-105.9-294.2,65.8
	c0,166.5,173.4,277.2,294.2,372.6C995.5,683.1,1173.8,566.7,1170.7,400.7z"/>
<path fill="#FFFFFF" d="M876.5,341.8c-76.7-161.2-295-105.9-294.2,65.8c0,166.5,173.4,277.2,294.2,372.6l0,0V341.8z"/>
<path fill="none" stroke="#00B7D3" stroke-width="2" stroke-miterlimit="10" d="M1170.7,400.7c-2.2-172.1-220.5-220.9-294.2-58.4
	c-76.7-161.2-295-105.9-294.2,65.8c0,166.5,173.4,277.2,294.2,372.6C995.5,683.1,1173.8,566.7,1170.7,400.7z"/>
</svg>
