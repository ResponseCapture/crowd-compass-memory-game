<svg xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" version="1.1" id="imgView" x="0px" y="0px" width="256px" height="256px" viewBox="0 0 430.117 430.118" style="enable-background:new 0 0 430.117 430.118;" xml:space="preserve">
<g>
  <path id="ShareThis" d="M151.804,215.059c0,1.475-0.336,2.856-0.423,4.326l154.111,77.03   c13.194-11.173,30.075-18.146,48.725-18.146c41.925,0.009,75.9,33.985,75.9,75.905c0,41.967-33.976,75.942-75.9,75.942   c-41.961,0-75.9-33.976-75.9-75.942c0-1.512,0.336-2.861,0.42-4.326l-154.111-77.035c-13.234,11.131-30.075,18.104-48.725,18.104   c-41.922,0-75.9-33.938-75.9-75.858c0-41.962,33.979-75.945,75.9-75.945c18.649,0,35.496,7.017,48.725,18.148l154.111-77.035   c-0.084-1.473-0.42-2.858-0.42-4.368c0-41.88,33.939-75.859,75.9-75.859c41.925,0,75.9,33.979,75.9,75.859   c0,41.959-33.976,75.945-75.9,75.945c-18.691,0-35.539-7.017-48.725-18.19l-154.111,77.077   C151.463,212.163,151.804,213.549,151.804,215.059z"></path>
</g>
</svg>