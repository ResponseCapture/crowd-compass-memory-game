<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 18.1.1, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
	 viewBox="0 0 300 35" enable-background="new 0 0 300 35" xml:space="preserve">
<g>
	<path fill="#283238" d="M1129.6,781.5c-2.5,0-3.6,1.4-4.2,2.3v0h0c0,0,0,0,0,0v-2h-4.7c0.1,1.3,0,14.1,0,14.1h4.7V788
		c0-0.4,0-0.8,0.2-1.1c0.3-0.8,1.1-1.7,2.4-1.7c1.7,0,2.4,1.3,2.4,3.2v7.5h4.7v-8.1C1134.9,783.5,1132.6,781.5,1129.6,781.5z"/>
	<path fill="#283238" d="M1115.7,775c-1.6,0-2.7,1.1-2.7,2.4c0,1.4,1,2.4,2.6,2.4h0c1.6,0,2.7-1.1,2.7-2.4
		C1118.3,776,1117.3,775,1115.7,775z"/>
	<rect x="1113.4" y="781.8" fill="#283238" width="4.7" height="14.1"/>
</g>
<g>
	<g>
		<g>
			<g>
				<g>
					<path fill="#FFFFFF" d="M37.3,10.5c5.3,0,9.6,4.1,9.9,9.4h3.9c-0.1-4-1-7.7-2.5-10.7c-3.2-1.6-7.1-2.5-11.3-2.5
						s-8.1,0.9-11.3,2.5c-1.5,3-2.4,6.7-2.5,10.7h3.9C27.7,14.6,32,10.5,37.3,10.5z"/>
					<path fill="#FFFFFF" d="M37.3,30.3c-5.3,0-9.6-4.1-9.9-9.4h-3.9c0.1,4,1,7.7,2.5,10.7c3.2,1.6,7.1,2.5,11.3,2.5
						s8.1-0.9,11.3-2.5c1.5-3,2.4-6.7,2.5-10.7h-3.9C46.9,26.1,42.6,30.3,37.3,30.3z"/>
				</g>
				<g>
					<path fill="#FFFFFF" d="M33.8,16.9L33.8,16.9L33.8,16.9l-3.5,10.5l10.5-3.5l0,0l0,0l3.5-10.5L33.8,16.9z M37.3,22.3
						c-1,0-1.9-0.8-1.9-1.9c0-1,0.8-1.9,1.9-1.9c1,0,1.9,0.8,1.9,1.9C39.2,21.4,38.4,22.3,37.3,22.3z"/>
				</g>
			</g>
			<g>
				<path fill="#FFFFFF" d="M74.1,22.5c-1,3.9-4.3,6.4-8.3,6.4c-5.1,0-8.6-4.1-8.6-8.5c0-4.2,3.2-8.5,8.6-8.5c5.1,0,7.9,4,8.3,6.5
					h-4.4c-0.5-1.2-1.7-2.9-4-2.9c-2.8,0-4.4,2.5-4.4,4.8c0,2.5,1.7,4.9,4.4,4.9c2.6,0,3.7-2.2,3.9-2.8H74.1z"/>
				<path fill="#FFFFFF" d="M75.5,16.4H79v1.3h0c0.3-0.6,1-1.7,3.1-1.7v3.7c-1.7,0-2.9,0.4-2.9,2.3v6.8h-3.7V16.4z"/>
				<path fill="#FFFFFF" d="M88.7,16c4.5,0,6.6,3.5,6.6,6.5c0,3-2.1,6.5-6.6,6.5c-4.5,0-6.6-3.5-6.6-6.5C82.1,19.5,84.3,16,88.7,16
					 M88.7,25.6c1.6,0,2.9-1.3,2.9-3.1c0-1.8-1.4-3.1-2.9-3.1c-1.6,0-2.9,1.3-2.9,3.1C85.8,24.3,87.1,25.6,88.7,25.6"/>
				<polygon fill="#FFFFFF" points="98.8,16.4 100.7,24 100.7,24 102.7,16.4 105.8,16.4 107.9,24 107.9,24 109.7,16.4 113.5,16.4 
					109.8,28.7 106.4,28.7 104.3,20.7 104.2,20.7 102.2,28.7 98.8,28.7 95,16.4 				"/>
				<path fill="#FFFFFF" d="M126.7,28.7h-3.5v-1.3h0c-0.3,0.5-1.2,1.7-3.7,1.7c-3.7,0-6.2-2.9-6.2-6.6c0-4.2,3-6.5,6.1-6.5
					c2.2,0,3.2,1.1,3.6,1.5v-5.1h3.7V28.7z M120.1,25.6c2.3,0,3.1-1.9,3.1-3.2c0-1.5-1.1-3.1-3.1-3.1c-2.1,0-3.1,1.7-3.1,3.1
					C117,24.4,118.4,25.6,120.1,25.6"/>
				<path fill="#FFFFFF" d="M144.7,22.5c-1,3.9-4.3,6.4-8.3,6.4c-5.1,0-8.6-4.1-8.6-8.5c0-4.2,3.2-8.5,8.6-8.5c5.1,0,7.9,4,8.3,6.5
					h-4.4c-0.5-1.2-1.7-2.9-4-2.9c-2.8,0-4.4,2.5-4.4,4.8c0,2.5,1.7,4.9,4.4,4.9c2.6,0,3.7-2.2,3.9-2.8H144.7z"/>
				<path fill="#FFFFFF" d="M152.2,16c4.5,0,6.6,3.5,6.6,6.5c0,3-2.1,6.5-6.6,6.5c-4.5,0-6.6-3.5-6.6-6.5
					C145.6,19.5,147.8,16,152.2,16 M152.2,25.6c1.6,0,2.9-1.3,2.9-3.1c0-1.8-1.4-3.1-2.9-3.1c-1.6,0-2.9,1.3-2.9,3.1
					C149.3,24.3,150.6,25.6,152.2,25.6"/>
				<path fill="#FFFFFF" d="M159.8,16.4h3.4v1.3h0c0.3-0.5,1.1-1.7,3.4-1.7c1.1,0,2.6,0.4,3.5,2.2c0.8-1.2,2-2.2,3.9-2.2
					c0.9,0,2.2,0.2,3.2,1.2c1.2,1.2,1.3,2,1.3,4.8v6.7H175v-6.5c0-1,0-2.7-1.9-2.7c-2,0-2,1.9-2,2.5v6.7h-3.7V22
					c0-0.7,0-2.6-1.8-2.6c-2.1,0-2.1,2-2.1,2.7v6.5h-3.7V16.4z"/>
				<path fill="#FFFFFF" d="M179.9,16.4h3.5v1.4h0h0c0.7-0.9,2-1.8,3.8-1.8c4.4,0,6,3.8,6,6.7c0,3.5-2.5,6.4-6,6.4
					c-2.2,0-3.3-1.1-3.7-1.5v5.2h-3.7V16.4z M189.6,22.5c0-1.5-1.1-3.1-3.1-3.1c-2,0-3.1,1.7-3.1,3.1c0,1.5,1.2,3.1,3.1,3.1
					C188.4,25.6,189.6,24.1,189.6,22.5"/>
				<path fill="#FFFFFF" d="M207.2,28.7h-3.7v-1.3h0c-0.6,1.2-2.1,1.7-3.6,1.7c-3.9,0-6.2-3.1-6.2-6.6c0-4,2.9-6.6,6.2-6.6
					c2,0,3.1,1,3.6,1.7h0v-1.3h3.7V28.7z M200.5,25.6c2.3,0,3.1-1.9,3.1-3.1c0-1.5-1-3.1-3.1-3.1c-2.1,0-3,1.8-3,3.2
					C197.4,23.7,198.3,25.6,200.5,25.6"/>
				<path fill="#FFFFFF" d="M214.3,19.8c0-0.3-0.1-0.9-1.2-0.9c-0.8,0-1,0.5-1,0.8c0,0.7,0.9,1,1.9,1.3c2.1,0.6,4.3,1.2,4.3,3.9
					c0,2.6-2.3,4.2-5,4.2c-1.9,0-4.7-0.8-5-4.1h3.7c0.2,1.1,1.2,1.1,1.4,1.1c0.6,0,1.3-0.4,1.3-1c0-1-0.9-1.1-3.3-2
					c-1.6-0.5-2.9-1.6-2.9-3.2c0-2.4,2.2-4.1,4.8-4.1c1.6,0,4.4,0.6,4.7,3.9H214.3z"/>
				<path fill="#FFFFFF" d="M224.7,19.8c0-0.3-0.1-0.9-1.2-0.9c-0.8,0-1,0.5-1,0.8c0,0.7,0.9,1,1.9,1.3c2.1,0.6,4.3,1.2,4.3,3.9
					c0,2.6-2.3,4.2-5,4.2c-1.9,0-4.7-0.8-5-4.1h3.7c0.2,1.1,1.2,1.1,1.4,1.1c0.6,0,1.3-0.4,1.3-1c0-1-0.9-1.1-3.3-2
					c-1.6-0.5-2.9-1.6-2.9-3.2c0-2.4,2.2-4.1,4.8-4.1c1.6,0,4.4,0.6,4.7,3.9H224.7z"/>
			</g>
		</g>
	</g>
	<g>
		<g>
			<g>
				<path fill="#FFFFFF" d="M235.7,28.6v-7.7h0.9v3c0.2-0.3,0.5-0.6,0.8-0.7c0.3-0.2,0.7-0.3,1.1-0.3c0.4,0,0.7,0.1,1,0.2
					c0.3,0.1,0.6,0.3,0.8,0.6c0.2,0.3,0.4,0.6,0.5,0.9c0.1,0.4,0.2,0.8,0.2,1.2c0,0.5-0.1,0.9-0.2,1.2c-0.1,0.4-0.3,0.7-0.5,0.9
					c-0.2,0.3-0.5,0.4-0.8,0.6c-0.3,0.1-0.6,0.2-1,0.2c-0.4,0-0.8-0.1-1.1-0.3c-0.3-0.2-0.6-0.4-0.8-0.7v0.8H235.7z M236.5,27.1
					c0.2,0.2,0.4,0.5,0.7,0.6c0.3,0.2,0.6,0.3,1,0.3c0.3,0,0.5-0.1,0.8-0.2c0.2-0.1,0.4-0.3,0.6-0.5c0.2-0.2,0.3-0.4,0.4-0.7
					c0.1-0.3,0.1-0.5,0.1-0.9c0-0.3,0-0.6-0.1-0.9c-0.1-0.3-0.2-0.5-0.4-0.7c-0.2-0.2-0.3-0.3-0.6-0.5c-0.2-0.1-0.5-0.2-0.8-0.2
					c-0.3,0-0.7,0.1-1,0.3c-0.3,0.2-0.5,0.4-0.7,0.6V27.1z"/>
				<path fill="#FFFFFF" d="M242.3,30c0.1,0,0.1,0.1,0.2,0.1c0.1,0,0.2,0,0.2,0c0.2,0,0.4,0,0.5-0.1c0.1-0.1,0.2-0.2,0.3-0.5
					l0.4-0.8l-2.3-5.7h0.9l1.9,4.6l1.9-4.6h1l-2.8,6.7c-0.2,0.4-0.4,0.7-0.7,0.9c-0.3,0.2-0.6,0.3-1,0.3c-0.1,0-0.2,0-0.3,0
					c-0.1,0-0.2,0-0.3-0.1L242.3,30z"/>
				<path fill="#FFFFFF" d="M254.8,28.7c-0.6,0-1.1-0.1-1.6-0.3c-0.5-0.2-0.9-0.5-1.3-0.8c-0.4-0.4-0.6-0.8-0.8-1.3
					c-0.2-0.5-0.3-1-0.3-1.6c0-0.6,0.1-1.1,0.3-1.6c0.2-0.5,0.5-0.9,0.8-1.3c0.4-0.4,0.8-0.6,1.3-0.8c0.5-0.2,1-0.3,1.6-0.3
					c0.3,0,0.7,0,0.9,0.1c0.3,0.1,0.6,0.2,0.8,0.3c0.2,0.1,0.5,0.3,0.7,0.5c0.2,0.2,0.4,0.4,0.5,0.6l-0.8,0.5
					c-0.2-0.3-0.5-0.6-0.9-0.8c-0.4-0.2-0.8-0.3-1.2-0.3c-0.4,0-0.8,0.1-1.2,0.2c-0.4,0.2-0.7,0.4-0.9,0.6c-0.3,0.3-0.5,0.6-0.6,1
					c-0.2,0.4-0.2,0.8-0.2,1.3c0,0.5,0.1,0.9,0.2,1.3c0.2,0.4,0.4,0.7,0.6,1c0.3,0.3,0.6,0.5,0.9,0.6c0.4,0.2,0.8,0.2,1.2,0.2
					c0.4,0,0.8-0.1,1.2-0.3c0.4-0.2,0.7-0.5,0.9-0.8l0.8,0.5c-0.3,0.4-0.7,0.8-1.2,1.1C256.1,28.6,255.5,28.7,254.8,28.7z"/>
				<path fill="#FFFFFF" d="M260.5,28.6l-2.3-5.6h0.9l1.9,4.6l1.9-4.6h1l-2.3,5.6H260.5z"/>
				<path fill="#FFFFFF" d="M267,28.7c-0.4,0-0.8-0.1-1.1-0.2c-0.3-0.1-0.6-0.3-0.9-0.6c-0.3-0.3-0.4-0.6-0.6-0.9
					c-0.1-0.4-0.2-0.8-0.2-1.2c0-0.4,0.1-0.8,0.2-1.1c0.1-0.4,0.3-0.7,0.6-0.9c0.2-0.3,0.5-0.5,0.9-0.6c0.3-0.2,0.7-0.2,1.1-0.2
					c0.4,0,0.8,0.1,1.1,0.2c0.3,0.2,0.6,0.4,0.8,0.6c0.2,0.3,0.4,0.6,0.5,1c0.1,0.4,0.2,0.8,0.2,1.2v0.2h-4.5c0,0.3,0.1,0.5,0.2,0.7
					c0.1,0.2,0.2,0.4,0.4,0.6c0.2,0.2,0.4,0.3,0.6,0.4c0.2,0.1,0.5,0.2,0.8,0.2c0.3,0,0.6-0.1,0.9-0.2c0.3-0.1,0.6-0.3,0.8-0.5
					l0.4,0.6c-0.3,0.3-0.6,0.5-1,0.6C267.9,28.7,267.5,28.7,267,28.7z M268.8,25.5c0-0.2,0-0.4-0.1-0.6c-0.1-0.2-0.2-0.4-0.3-0.6
					c-0.2-0.2-0.3-0.3-0.6-0.4c-0.2-0.1-0.5-0.2-0.8-0.2c-0.3,0-0.6,0.1-0.8,0.2c-0.2,0.1-0.4,0.3-0.6,0.4c-0.2,0.2-0.3,0.4-0.3,0.6
					c-0.1,0.2-0.1,0.4-0.1,0.7H268.8z"/>
				<path fill="#FFFFFF" d="M274.6,28.6v-3.7c0-0.5-0.1-0.8-0.3-1c-0.2-0.2-0.5-0.3-0.9-0.3c-0.2,0-0.3,0-0.5,0.1
					c-0.2,0-0.3,0.1-0.5,0.2c-0.1,0.1-0.3,0.2-0.4,0.3c-0.1,0.1-0.2,0.2-0.3,0.3v4.1h-0.9V23h0.9v0.8c0.1-0.1,0.2-0.2,0.4-0.3
					c0.1-0.1,0.3-0.2,0.5-0.3c0.2-0.1,0.4-0.2,0.6-0.2c0.2-0.1,0.4-0.1,0.6-0.1c1.2,0,1.8,0.6,1.8,1.8v3.9H274.6z"/>
				<path fill="#FFFFFF" d="M278.5,28.7c-0.4,0-0.7-0.1-0.9-0.3c-0.2-0.2-0.3-0.5-0.3-1v-3.7h-0.9V23h0.9v-1.5h0.9V23h1.1v0.8h-1.1
					v3.5c0,0.2,0,0.4,0.1,0.5c0.1,0.1,0.2,0.2,0.4,0.2c0.1,0,0.2,0,0.3-0.1c0.1,0,0.2-0.1,0.2-0.2l0.3,0.6c-0.1,0.1-0.2,0.2-0.4,0.3
					C279,28.7,278.8,28.7,278.5,28.7z"/>
			</g>
		</g>
	</g>
</g>
</svg>
